//day3 is for rising_falling_edge_detector
